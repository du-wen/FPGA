module spi_ctrl(
    input   wire            sclk,//50M
    input   wire            rst_n,
    input   wire            work_en,//�������ò�����ʹ��
    output  reg             conf_end,//������ɱ�־
    output  wire            spi_clk,//50-60mhz
    output  wire            spi_sdi,
    output  wire            spi_csn,
    input   wire            spi_sdo//������ܽŲ����б��
);

parameter       IDLE = 5'b0_0001;
parameter       WAIT = 5'b0_0010;
parameter       R_MEM= 5'b0_0100;
parameter       W_REG= 5'b0_1000;
parameter       STOP = 5'b1_0000;
 
parameter       H_DIV_CYC   =   5'd25-1;//��Ƶ,���ڲ���1Mʱ��

reg     [4:0]   state;//״̬���ļĴ������������뷽ʽ���ö�����
reg     [4:0]   div_cnt;
reg             clk_p = 1'b0;
wire            clk_n;
reg             pose_flag;//���ڱ�־������
reg  [3:0]      wait_cnt;
reg  [3:0]      shift_cnt;
reg  [4:0]      r_addr;
wire [15:0]     r_data;
wire            wren;
reg  [15:0]     shift_buf;//��λ�Ĵ��������ڻ���ram��������ݣ���R_MEM״̬����ɸ�ֵ
reg            data_end;
reg             sdi;//spi������Ĵ���
reg             csn;
reg             tck;//����D��������ʱһ�ģ�ʹʱ�����������sdi���Ķ���

//��Ƶ������
always @(posedge sclk or negedge rst_n)
begin
  if (rst_n == 1'b0)
    div_cnt <= 5'd0;
  else if(div_cnt == H_DIV_CYC)
    div_cnt <= 5'd0;
  else
    div_cnt <= div_cnt + 1'b1;
end
//��Ƶʱ�Ӳ��������Ĵ����Ĵ���ʱ�ӣ�Ҳ���ǲ���д��always�Ĵ����б���(��׼ȷ)
always @(posedge sclk or negedge rst_n)
begin
  if(rst_n == 1'b0)
    clk_p <= 1'b0;
  else if(div_cnt == H_DIV_CYC)
    clk_p <= ~clk_p;
end

assign clk_n = ~clk_p;//������Ϊ�˴ﵽ���Ķ����Ŀ��

always @(posedge sclk or negedge rst_n)
begin
  if(rst_n == 1'b0)
    pose_flag <= 1'b0;
  else if(clk_p == 1'b0 && div_cnt == H_DIV_CYC)
    pose_flag <= 1'b1;         //clk_p���������ص�ʱ��pose_flag����,pose_flag����Ϊ1mhz����ʱ��Ϊ20ns������
  else  pose_flag <= 1'b0;
end

always @(posedge sclk or negedge rst_n)
  if(rst_n == 1'b0)
    wait_cnt <= 4'd0;
  else if (state == WAIT && pose_flag == 1'b1)
    wait_cnt <= wait_cnt + 1'b1;
  else if(state != WAIT)
    wait_cnt <= 4'd0;

//fsm���˴�������ʽ״̬��
always @(posedge sclk or negedge rst_n)
  if(rst_n == 1'b0)
    state <= IDLE;
  else case(state)
    IDLE: if(work_en == 1'b1)
            state <= WAIT;
    WAIT: if(wait_cnt[3] == 1'b1)
            state <= R_MEM;
    R_MEM: state <= W_REG;
    W_REG:if((shift_cnt == 4'd15) && (pose_flag == 1'b1 )&& (data_end != 1'b1))
            state <= WAIT;
          else if((shift_cnt == 4'd15) && (pose_flag == 1'b1 )&& (data_end == 1'b1))
            state <= STOP;
    STOP: state <= STOP;
    default: state <= IDLE;
  endcase

always @(posedge sclk or negedge rst_n)
  if(rst_n == 1'b0)
    shift_cnt <= 4'd0;
  else if(state == W_REG && pose_flag == 1'b1)
    shift_cnt <= shift_cnt + 1'b1;
  else if(state != W_REG)
    shift_cnt <= 4'd0;

//��mem�ĵ�ַ�Ĳ�������R_MEMʱ�򾭹�D��������ֵ����W_REGʵ�ֵ�ַ��1
always @(posedge sclk or negedge rst_n)
  if(rst_n == 1'b0)
    r_addr <=  4'd0;
  else if(state == R_MEM)
    r_addr <= r_addr + 1'b1;

//data_end���һ����Ҫ��λ����
always @(posedge sclk or negedge rst_n)
  if(rst_n == 1'b0)
    data_end <= 5'd0;
  else if(state == R_MEM && (&r_addr) == 1'b1)//��Ч��state == R_MEM && r_addr == 5'd31
    data_end <= 1'b1;


assign wren = 1'b0;  

always @(posedge sclk or negedge rst_n)
   if(rst_n == 1'b0)
     shift_buf <= 16'd0;
   else if(state == R_MEM)
     shift_buf <= r_data;//R_MEM״̬�£����ݻ������
   else if(state == W_REG && pose_flag == 1'b1)
     shift_buf <= {shift_buf[14:0],1'b1};//W_REG��pose_flagΪ1ʱ����������һλ���Ƶ�sdi��ȥ���൱�ڲ�ת����

//�������
always @(posedge sclk or negedge rst_n)
  if(rst_n == 1'b0)
    sdi <= 1'b0;
  else if(state == W_REG)//����state == W_REG && pose_flag == 1'b1,��sclkͬ������������pose_flagͬ���������Ӻ�sclk��������pose_flag��ʹ�����һλ���ݾ����ٴ���STOP״̬��
    sdi <= shift_buf[15];
  else if(state != W_REG)
    sdi <= 1'b0;
    
//cs�Ĳ�������sdi����
always @(posedge sclk or negedge rst_n)
  if(rst_n == 1'b0)
    csn <= 1'b1;//csnΪ0ʱ��ѡͨ
  else if(state == W_REG)
    csn <= 1'b0;
  else 
    csn <= 1'b1;  

//�������������Ķ����ʱ��
always @(posedge sclk or negedge rst_n)
  if(rst_n == 1'b0)
    tck <= 1'b0;
  else if(state == W_REG)//state����־��
    tck <= clk_n;
  else
    tck <= 1'b0;

assign spi_clk = tck;
assign spi_csn = csn;
assign spi_sdi = sdi;

always @(posedge sclk or negedge rst_n)
  if(rst_n == 1'b0)
    conf_end <= 1'b0;
  else if(state == STOP)
    conf_end <= 1'b1;
    
//��ram��rom�ã����ǲ��������д������ֻ�ǲ��ϵĴ�ram�ж�����
ram_16_32_sr	ram_16_32_sr_inst (
	.address ( r_addr ),//����ַ
	.clock ( sclk ),
	.data ( 16'd0 ),//д����
	.wren ( wren ),//дʹ�ܸ���Ч����ʹ�ܵ���Ч
	.q ( r_data )//������
	);
    
//ȫ����sclk��Ϊʱ�ӣ����ü�����������clk_pʱ�ӣ�sclk��ϵͳʱ�ӣ��᲼�ֵ�ȫ��ʱ�����磬clk_p��Ϊ�����ߣ�������ܴ��ʱ��ƫб��skew������Ӱ�����ǵĽ���ʱ�������ʱ�䡣��ˣ�������sclk��Ϊͬ��ʱ�ӡ� 
endmodule